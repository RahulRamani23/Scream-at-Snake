module game_overlay(
    output [2699:0] OUT, 
    input is_high_score,
    input is_win,
    input clock
);

    wire [699:0] game_over_text_wire, motivation_text_wire;
    wire [499:0] high_score_winner_wire;
    wire [199:0] line_break;

    assign line_break = 300'd0;

    game_over_text game_over (
        .OUT(game_over_text_wire)
    );

    high_score_winner_text high_score_winner (
        .OUT(high_score_winner_wire),
        .is_high_score(is_high_score),
        .is_win(is_win),
        .clock(clock)
    );

    motivation_text motivation (
        .OUT(motivation_text_wire),
        .is_high_score(is_high_score),
        .is_win(is_win),
        .clock(clock)
    );

    assign OUT = {high_score_winner_wire, line_break, motivation_text_wire, line_break, game_over_text_wire};

    
endmodule


module game_over_text(
    output [699:0] OUT
);
	// Changed this text to R.I.P.
    assign OUT[99:0] 	= 100'b0000000000000000000000011111111100000000000000011111111110000000000011111111100000000000000000000000;
    assign OUT[199:100] = 100'b0000000000000000000000100000001100000000000000000001100000000000000100000001100000000000000000000000;
    assign OUT[299:200] = 100'b0000000000000000000000100000001100000000000000000001100000000000000010000001100000000000000000000000;
    assign OUT[399:300] = 100'b0000000000000000000000011111111100000000000000000001100000000000000001111111100000000000000000000000;
    assign OUT[499:400] = 100'b0000000000000000000000000000001100000000000000000001100000000000000000000101100000000000000000000000;
    assign OUT[599:500] = 100'b0000000000000000110000000000001100000011000000000001100000000011000000001001100000000000000000000000;
    assign OUT[699:600] = 100'b0000000000000000110000000000001100000011000000011111111110000011000000110001100000000000000000000000;





endmodule

module high_score_winner_text(
    output reg [499:0] OUT,
    input is_high_score,
    input is_win,
    input clock
);

    wire clear = 500'd0;

    always@(*)
    begin
        if(is_win)
            begin
                OUT[99:0] 		= 100'b0000000000000000000000000000000000000111101111010011010011010100010000000000000000000000000000000000;
                OUT[199:100] 	= 100'b0000000000000000000000000000000000001000100001010101010101010100010000000000000000000000000000000000;
                OUT[299:200] 	= 100'b0000000000000000000000000000000000000111100011011001011001010101010000000000000000000000000000000000;
                OUT[399:300] 	= 100'b0000000000000000000000000000000000000100100001010001010001010110110000000000000000000000000000000000;
                OUT[499:400] 	= 100'b0000000000000000000000000000000000001000101111010001010001010100010000000000000000000000000000000000;
            end
        else if(is_high_score)
            begin
                OUT[99:0] 		= 100'b0000000000000000000000011110001111001111000111000111000010001011110001001000100000000000000000000000;
                OUT[199:100] 	= 100'b0000000000000000000000000010010001010000101000100000100010001000001001001000100000000000000000000000;
                OUT[299:200] 	= 100'b0000000000000000000000001110001001010000100000100011000011111010001001001111100000000000000000000000;
                OUT[399:300] 	= 100'b0000000000000000000000000010010001010000101000100100000010001010001001001000100000000000000000000000;
                OUT[499:400] 	= 100'b0000000000000000000000011110100001001111000111000111100010001001110001001000100000000000000000000000;
            end
			else
				OUT = clear;
    end
endmodule


module motivation_text(
    output reg [699:0] OUT,
    input is_high_score,
    input is_win,
    input clock
);
    wire [1:0] random_3;

    random generator(
        .clock(clock),
        .max_number(2'b10),
        .num_out(random_3)
    );

    wire [699:0] motivation_1, motivation_2, motivation_3;
    wire [699:0] success_1, success_2, success_3;
    wire [699:0] win;

    // Changed to GO HOME
    assign motivation_1[99:0] 	= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign motivation_1[199:100] = 100'b0000000000000000000000011110000100010000011100001001000000000001110000111100000000000000000000000000;
    assign motivation_1[299:200] = 100'b0000000000000000000000000010000110110000100010001001000000000010001000000100000000000000000000000000;
    assign motivation_1[399:300] = 100'b0000000000000000000000001110000101010000100010001111000000000010001000110100000000000000000000000000;
    assign motivation_1[499:400] = 100'b0000000000000000000000000010000100010000100010001001000000000010001000100100000000000000000000000000;
    assign motivation_1[599:500] = 100'b0000000000000000000000011110000100010000011100001001000000000001110000111100000000000000000000000000;
    assign motivation_1[699:600] = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // Changed to YIKES
    assign motivation_2[99:0] 	= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign motivation_2[199:100] = 100'b0000000000000000000000000000011100000001111000010010000010000001000100000000000000000000000000000000;
    assign motivation_2[299:200] = 100'b0000000000000000000000000000000010000000001000001010000010000000101000000000000000000000000000000000;
    assign motivation_2[399:300] = 100'b0000000000000000000000000000011100000000111000000110000010000000010000000000000000000000000000000000;
    assign motivation_2[499:400] = 100'b0000000000000000000000000000010000000000001000001010000010000000010000000000000000000000000000000000;
    assign motivation_2[599:500] = 100'b0000000000000000000000000000001110000001111000010010000010000000010000000000000000000000000000000000;
    assign motivation_2[699:600] = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // changed toPress F!
    assign motivation_3[99:0] 	= 100'b0000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign motivation_3[199:100] = 100'b0000000000001111100000011111111111110000000000000000000000000000000000000000111111000000000000000000;
    assign motivation_3[299:200] = 100'b0000000000000111000000000000000000110000000000000000011000110001110000111100110001100000000000000000;
    assign motivation_3[399:300] = 100'b0000000000000111000000000000011111110000000000000000000100001001001001001100011111100000000000000000;
    assign motivation_3[499:400] = 100'b0000000000000000000000000000000000110000000000000000001000010000111000001100000001100000000000000000;
    assign motivation_3[599:500] = 100'b0000000000000111000000000000000000110000000000000000010000100000001000001100000001100000000000000000;
    assign motivation_3[699:600] = 100'b0000000000000111000000000000000000110000000000000000001100011001110000001100000001100000000000000000;

    // changed to 1001001 (this a reference to the big bang theory as an easter egg)
    assign success_1[99:0] 	= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign success_1[199:100] = 100'b0000000000000011000000000111000000000111000000000110000000001110000000001110000000001100000000000000;
    assign success_1[299:200] = 100'b0000000000000011000000001000100000001000100000000110000000010001000000010001000000001100000000000000;
    assign success_1[399:300] = 100'b0000000000000011000000010000010000010000010000000110000000100000100000100000100000001100000000000000;
    assign success_1[499:400] = 100'b0000000000000011000000001000100000001000100000000110000000010001000000010001000000001100000000000000;
    assign success_1[599:500] = 100'b0000000000000011000000000111000000000111000000000110000000001110000000001110000000001100000000000000;
    assign success_1[699:600] = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // Changed to Brian Approves!
    assign success_2[99:0] 	= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign success_2[199:100] = 100'b0000001100000111000011110000100010000011100001110001110011100111000001000100011100010001110001110000;
    assign success_2[299:200] = 100'b0000001100000000100000010000100010000100010010010010010100101000100001001100100010010010010010010000;
    assign success_2[399:300] = 100'b0000001100000111100001110000010100000100010001110011110111101110100001010100111010010001110001110000;
    assign success_2[499:400] = 100'b0000000000000100000000010000010100000100010001010000010000101000100001100100100010010001010010010000;
    assign success_2[599:500] = 100'b0000001100000011100011110000001000000011100010010000010000101000100001000100100010010010010001110000;
    assign success_2[699:600] = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // Changed to DANK!!
    assign success_3[99:0] 	= 100'd0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign success_3[199:100] = 100'b0000000000000000000000000000110011000000010100000100010000001110000000011100000000000000000000000000;
    assign success_3[299:200] = 100'b0000000000000000000000000000110011000000010100000100110000010001000000100100000000000000000000000000;
    assign success_3[399:300] = 100'b0000000000000000000000000000110011000000001100000101010000011101000000100100000000000000000000000000;
    assign success_3[499:400] = 100'b0000000000000000000000000000000000000000010100000110010000010001000000100100000000000000000000000000;
    assign success_3[599:500] = 100'b0000000000000000000000000000110011000000010100000100010000010001000000011100000000000000000000000000;
    assign success_3[699:600] = 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // Unbelievable
    assign win[99:0] 	= 100'd0;
    assign win[199:100] = 100'b0000000000000000000000100000001000001000000000000000000101000000000010000001001000000000000000000000;
    assign win[299:200] = 100'b0000000000000000000000100000001000001000000000000000000001000000000010000001001000000000000000000000;
    assign win[399:300] = 100'b0000000000000000000000100111001001101001111000000011100101011100011010011101001000000000000000000000;
    assign win[499:400] = 100'b0000000000000000000000100111101010011011110010001011110101011110100110100101001000000000000000000000;
    assign win[599:500] = 100'b0000000000000000000000000000101010001010001001010000010101000010100010100101001000000000000000000000;
    assign win[699:600] = 100'b0000000000000000000000100111001001111011110000100011100101011100011110100100110000000000000000000000;

    always @(*)
    begin
        if (is_win == 1'b1)
            OUT = win;
        else if (is_high_score == 1'b1)
            case(random_3[1:0])
                2'b00: OUT = success_1;
                2'b01: OUT = success_2;
                2'b10: OUT = success_3;
					 default: OUT = success_1;
            endcase
        else
            case(random_3[1:0])
                2'b00: OUT = motivation_1;
                2'b01: OUT = motivation_2;
                2'b10: OUT = motivation_3;
					default: OUT = motivation_1;
            endcase
    end
endmodule
